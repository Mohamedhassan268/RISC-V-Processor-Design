module Mux2_32 (
    input  [31:0] a,
    input  [31:0] b,
    input         sel,
    output [31:0] y
);

    // 👉 your assign line will go here

endmodule
