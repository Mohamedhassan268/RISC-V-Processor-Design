module Adder32 (
    input  [31:0] a,
    input  [31:0] b,
    output [31:0] y
);

    // ?? YOUR LINE GOES HERE

endmodule

